//////////////////////////////////////////////////////////////////////////////////
// Company:         UW
// Engineer:        Henry Wysong-Grass
// 
// Create Date:     2026-02-12
// Design Name:     SPART (Special Purpose Asynchronous Receiver/Transmitter)
// Module Name:     spart 
//
// Revision: 
// Revision 1.00 - Dummy implementation
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


module spart(
    input clk,
    input rst,
    input iocs,
    input iorw,
    output rda,
    output tbr,
    input [1:0] ioaddr,
    inout [7:0] databus,
    output txd,
    input rxd
    );





endmodule
