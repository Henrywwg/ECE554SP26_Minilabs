module bus_interface(
    
);



endmodule