// Matrix-vector multiplier

module matvec_mult (
    input logic clk,
    input logic rst_n,
    input logic 
);


endmodule